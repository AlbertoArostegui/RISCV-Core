`define PC_INITIAL 32'h00000000

`define OPCODE_RTYPE    7'b0110011
`define OPCODE_STORE    7'b0100011
`define OPCODE_LOAD     7'b0000011
`define OPCODE_JUMP     7'b1101111
`define OPCODE_BRANCH   7'b1100011
