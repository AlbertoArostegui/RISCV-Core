module imemory (
    input clk,
    input [31:0] mem_addr,
    output [31:0] inst_out
);

    reg [31:0] ROM [0:1023];

    initial begin
        ROM[0] = 32'b0000000_00010_00011_000_00001_0110011; //add r1, r2, r3
        ROM[1] = 32'b0000000_00010_00001_000_00001_0110011; //add r1, r2, r1
        ROM[2] = 32'b00000000_00000000_00000000_00000011;
        ROM[3] = 32'b00000000_00000000_00000000_00000001;
        ROM[4] = 32'b00000000_00000000_00000000_00000001;
        ROM[5] = 32'b00000000_00000000_00000000_00000001;
        ROM[6] = 32'b00000000_00000000_00000000_00000011;
        ROM[7] = 32'b00000000_00000000_00000000_00000111;
        ROM[8] = 32'b00000000_00000000_00000000_00001111;
        ROM[9] = 32'b00000000_00000000_00000000_00000011;
        ROM[10] = 32'b00000000_00000000_00000000_00000011;
        ROM[11] = 32'b00000000_00000000_00000000_00000011;
        ROM[12] = 32'b00000000_00000000_00000000_00000011;
        ROM[13] = 32'b00000000_00000000_00000000_00000011;
        ROM[14] = 32'b00000000_00000000_00000000_00000011;
        ROM[15] = 32'b00000000_00000000_00000000_00000011;
    end

    assign inst_out = ROM[mem_addr];

endmodule
