`define PC_INITIAL 32'h0
