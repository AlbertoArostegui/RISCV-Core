module imemory (
    input clk,
    input [31:0] mem_addr,
    output [31:0] inst_out
);

    reg [31:0] ROM [0:1023];

    initial begin
        ROM[0] = 32'b0000000_00010_00011_000_00001_0110011; //add r1, r2, r3
        ROM[1] = 32'b0000000_00110_00101_000_00100_0110011; //add r4, r5, r6
        ROM[2] = 32'b0000000_00010_00011_000_00001_0110011;
        ROM[3] = 32'b0000000_00010_00011_000_00001_0110011;
        ROM[4] = 32'b0000000_00010_00011_000_00001_0110011;
        ROM[5] = 32'b0000000_00010_00011_000_00001_0110011;
        ROM[6] = 32'b0000000_00010_00011_000_00001_0110011;
        ROM[7] = 32'b0000000_00010_00011_000_00001_0110011;
        ROM[8] = 32'b0000000_00010_00011_000_00001_0110011;
        ROM[9] = 32'b0000000_00010_00011_000_00001_0110011;
   end

    assign inst_out = ROM[mem_addr];

endmodule
