module reorder_buffer(
    input clk,
    input reset,

);

endmodule
